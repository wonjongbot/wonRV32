module soc (
    input logic clk,
    input logic reset,
    output logic
